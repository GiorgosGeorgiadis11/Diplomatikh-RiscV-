LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY WORK;
USE WORK.TOOLBOX.ALL;

ENTITY SIZE_COMPARATOR IS

	PORT(
		A : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		B : IN  STD_LOGIC_VECTOR(31  DOWNTO 0);
		O : OUT STD_LOGIC
	    );
		 
END SIZE_COMPARATOR;

ARCHITECTURE STRUCTURAL OF SIZE_COMPARATOR IS
	SIGNAL A_EXTENDED : STD_LOGIC_VECTOR(32 DOWNTO 0);
	SIGNAL B_EXTENDED : STD_LOGIC_VECTOR(32 DOWNTO 0);
	SIGNAL SUB_RES : STD_LOGIC_VECTOR(32 DOWNTO 0);
    BEGIN
		A_EXTENDED <= '0' & A;
		B_EXTENDED <= '0' & B;
		Sub: EXE_ADDER_SUBBER --(A-B)
		PORT MAP(
				A  => A_EXTENDED,
				B  => B_EXTENDED,
				OP => '1',
				S  => SUB_RES
			);
		-- if A-B < 0 then SUB_RES(32) while be 1 else while be 0
		O <= NOT SUB_RES(32); -- if A>=B return 1 else return 0
END STRUCTURAL;
