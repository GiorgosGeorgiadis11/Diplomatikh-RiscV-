-- +===========================================================+
-- |		RISC-V RV32I(M) ISA IMPLEMENTATION  	           |
-- |===========================================================|
-- |student:    Georgios Georgiadis			                   |
-- |supervisor: Kavousianos Xrysovalantis			           |
-- |===========================================================|
-- |		UNIVERSITY OF IOANNINA - 2022      	               |
-- |  		     VCAS LABORATORY			                   |
-- +===========================================================+

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;	
USE IEEE.STD_LOGIC_MISC.ALL;

LIBRARY WORK;
USE WORK.TOOLBOX.ALL;

ENTITY EXE_MUL_DIV IS 

	PORT(
		MULTICYCLING : IN STD_LOGIC;
		A  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		B  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		OP : IN  STD_LOGIC_VECTOR(9  DOWNTO 0);
        CYCLE : IN  STD_LOGIC_VECTOR(4  DOWNTO 0);
        PREVPCS : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
        PREVPCC : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
        PREVRESULT : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        ISMULDIV : OUT STD_LOGIC;
        NEXTPCS : OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
        NEXTPCC : OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		NEXTRESULT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		RES  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
			
	    );

END EXE_MUL_DIV;

ARCHITECTURE STRUCTURAL OF EXE_MUL_DIV IS 
	-- MUL/DIV SIGS ----------------------------
	SIGNAL A_COMPLEMENT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL B_COMPLEMENT : STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL END_MULTICYCLING : STD_LOGIC;
	SIGNAL END_MULTICYCLING_DIV : STD_LOGIC;
	SIGNAL END_MULTICYCLING_MUL : STD_LOGIC;
	SIGNAL END_CYCLE :STD_LOGIC;

	SIGNAL NEXTPCSMUL : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NEXTPCSDIV : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NEXTRESULTMUL : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NEXTRESULTDIV : STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL DIV_COMPLEMENT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REM_COMPLEMENT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MUL_COMPLEMENT : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MULH_COMPLEMENT: STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL MUL_RES    : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MULH_RES   : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL DIV_RES    : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REM_RES    : STD_LOGIC_VECTOR(31 DOWNTO 0);

	SIGNAL RESZERO32 : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
	BEGIN
		
	--MULTICYCLING MUL/DIV
	END_MULTICYCLING_MUL <= AND_REDUCE(CYCLE(1 DOWNTO 0)); -- 4 CYCLES MULTIPLICATION
	--END_MULTICYCLING_MUL <= CYCLE(0); -- 2 CYCLES MULTIPLICATION
	END_MULTICYCLING_DIV <= AND_REDUCE(CYCLE(4 DOWNTO 0)); -- 32 CYCLES DIVISION
	--END_MULTICYCLING_DIV <= AND_REDUCE(CYCLE(3 DOWNTO 0)); -- 16 CYCLES DIVISION

	END_MULTICYCLING_CYCLE: MUX2X1_BIT
		PORT MAP(
				D0  => END_MULTICYCLING_MUL,
				D1  => END_MULTICYCLING_DIV,
				SEL => OP(6),
				O   => END_CYCLE
			);
	END_MULTICYCLING <= NOT (END_CYCLE AND OP(7));

	-- TWO_COMPLEMENT ---------------------------------
	ISMULDIV <= END_MULTICYCLING AND OP(7) AND MULTICYCLING;

	TWO_COMPLEMENT_BEFORE: TWOS_COMPLEMENT
		PORT MAP(
			A  => A,
			B  => B,
			SIGNA  => A(31),
			SIGNB  => B(31),
			BEFOREAFTER  => '0',
			OP  => OP(9 DOWNTO 8),
			ONEREGMANAGMENT => '0',
			RESULTA => A_COMPLEMENT,
			RESULTB => B_COMPLEMENT
		);

    
	--ONE CYCLE MUL ---------------------------------
	-- --i_MUL: BASIC_MUL
	-- --i_MUL: ARRAY_MUL
	-- i_MUL: RIPPLE_CARRY_MUL
	-- 	PORT MAP(
	-- 			A => A_COMPLEMENT,
    --             B => B_COMPLEMENT,
	-- 			MSBRESULT => MULH_COMPLEMENT,
	-- 			RESULT => MUL_COMPLEMENT
	-- 		);
	--MULTICYCLING MUL ---------------------------------
	i_MUL: MUL_MULTICYCLING
		PORT MAP(
				A => A_COMPLEMENT,
                B => B_COMPLEMENT,
				PREVPCS => PREVPCS,
                PREVPCC => PREVPCC,
                PREVRESULT => PREVRESULT,
                CYCLE => CYCLE,
                NEXTPCS => NEXTPCSMUL,
                NEXTPCC => NEXTPCC,
				NEXTRESULT => NEXTRESULTMUL,
				MSBRESULT => MULH_COMPLEMENT,
				RESULT => MUL_COMPLEMENT
			);
	TWO_COMPLEMENT_MUL_AFTER: TWOS_COMPLEMENT
		PORT MAP(
			A  => MUL_COMPLEMENT,
			B  => MULH_COMPLEMENT,
			SIGNA  => A(31),
			SIGNB  => B(31),
			BEFOREAFTER  => '1',
			OP  => OP(9 DOWNTO 8),
			ONEREGMANAGMENT => '1',
			RESULTA => MUL_RES,
			RESULTB => MULH_RES
		);
    
	-- ONE CYCLE DIV ---------------------------------
	-- --i_DIV: LONG_DIV
	-- --i_DIV: IMPROVE_LONG_DIV
	-- i_DIV: ARRAY_DIV
	-- 	PORT MAP(
	-- 		A => A_COMPLEMENT,
    --         B => B_COMPLEMENT,
	-- 		REMAINDER => REM_COMPLEMENT,
    --         RESULT => DIV_COMPLEMENT  
	-- 	);	
	-- MULTICYCLING DIV ---------------------------------
	i_DIV: DIV_MULTICYCLING
		PORT MAP(
			A => A_COMPLEMENT,
            B => B_COMPLEMENT,
            PREVPCS => PREVPCS,
            PREVRESULT => PREVRESULT,
            CYCLE => CYCLE,
            NEXTPCS => NEXTPCSDIV,
			NEXTRESULT => NEXTRESULTDIV,
            RESULT => DIV_COMPLEMENT,
            REMAINDER => REM_COMPLEMENT
            
		);
	TWO_COMPLEMENT_DIV_AFTER: TWOS_COMPLEMENT
		PORT MAP(
			A  => DIV_COMPLEMENT,
			B  => REM_COMPLEMENT,
			SIGNA  => A(31),
			SIGNB  => B(31),
			BEFOREAFTER  => '1',
			OP  => OP(9 DOWNTO 8),
			ONEREGMANAGMENT => '0',
			RESULTA => DIV_RES,
			RESULTB => REM_RES
		);
	
	NEXTPCS_MUX: MUX2X1
        GENERIC MAP( INSIZE => 32 )
        PORT    MAP( 
                D0  => NEXTPCSMUL,
                D1  => NEXTPCSDIV,
                SEL => OP(6),
                O   => NEXTPCS
                );
	NEXTRESULT_MUX: MUX2X1
		GENERIC MAP( INSIZE => 32 )
		PORT    MAP( 
				D0  => NEXTRESULTMUL,
				D1  => NEXTRESULTDIV,
				SEL => OP(6),
				O   => NEXTRESULT
				);
				
	ALU_MUX: MUX4X1
		GENERIC MAP( INSIZE => 32 )
		PORT    MAP( 
				D0  => MUL_RES,
				D1  => MULH_RES,
				D2  => DIV_RES,
				D3  => REM_RES,
				SEL => OP(6 DOWNTO 5),
				O   => RES
				);		
END STRUCTURAL;