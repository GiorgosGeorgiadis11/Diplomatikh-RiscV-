LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

LIBRARY WORK;
USE WORK.TOOLBOX.ALL;

ENTITY SIZE_COMPARATOR IS

	PORT(
		A : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		B : IN  STD_LOGIC_VECTOR(31  DOWNTO 0);
		O : OUT STD_LOGIC
	    );
		 
END SIZE_COMPARATOR;

ARCHITECTURE RTL OF SIZE_COMPARATOR IS

    BEGIN
        PROCESS(A,B)
        BEGIN
            IF A>=B THEN
                O<='1';
            ELSE
                O<='0';
            END IF;

        END PROCESS;


END RTL;
