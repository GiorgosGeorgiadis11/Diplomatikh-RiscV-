LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

LIBRARY WORK;
USE WORK.TOOLBOX.ALL;

ENTITY MUL IS

	PORT(
		  A : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		  B : IN  STD_LOGIC_VECTOR(31  DOWNTO 0);
		  RESULT  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	    );
		 
END MUL;

ARCHITECTURE STRUCTURAL OF MUL IS
    TYPE ARR4 IS ARRAY(0 TO 32) OF STD_LOGIC_VECTOR(4 DOWNTO 0);
    TYPE ARR31 IS ARRAY(0 TO 32) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
    TYPE ARR32 IS ARRAY(0 TO 32) OF STD_LOGIC_VECTOR(32 DOWNTO 0);
    SIGNAL SHAMT  : ARR4;
    SIGNAL MUXOUT : ARR31;
    SIGNAL OUTPUT : ARR31;
    SIGNAL OUTPUTEXTENDED : ARR32;
    SIGNAL FINALOUT : ARR32;
    SIGNAL RESZERO : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
    SIGNAL OPADD  : STD_LOGIC := '0';
    SIGNAL OPSFT  : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
  
	BEGIN
    MAIN: FOR I IN 0 TO 31 GENERATE
      CHECKONE :MUX2X1
        GENERIC MAP(INSIZE => 32)
          PORT MAP(
            D0 => RESZERO,
            D1 => B,
            SEL => A(I),
            O=> MUXOUT(I)
          );
          
      INITIALIZE: IF I = 0 GENERATE
        FINALOUT(I)<=(OTHERS=>'0');
        OUTPUT(I)<=MUXOUT(I);
        SHAMT(I)<="00001";
      END GENERATE INITIALIZE;
      
      SFT: IF I > 0 GENERATE
        SHAMT(I)<=std_logic_vector(unsigned(SHAMT(I-1)) + 1);
        SHIFTER :BARREL_SHIFTER
          PORT MAP(
            VALUE_A =>MUXOUT(I),
            SHAMT_B =>SHAMT(I-1),
            OPCODE =>OPSFT,
            RESULT =>OUTPUT(I)
          );
      END GENERATE SFT;   
      OUTPUTEXTENDED(I)<='0'&OUTPUT(I);
      OUTPUTADD :EXE_ADDER_SUBBER
        PORT MAP(
          A=>OUTPUTEXTENDED(I),
          B=>FINALOUT(I),
          OP=>OPADD,
          S=>FINALOUT(I+1)
        );
        
    END GENERATE MAIN;
    RESULT<=FINALOUT(32)(31 DOWNTO 0);
        
END STRUCTURAL;
